module prencoder_32_5(in,y);
input[31:0] in;
output reg[4:0] y;

always@*
begin
casex(in)
32'b00000000000000000000000000000001:y=5'b00000;
32'b0000000000000000000000000000001x:y=5'b00001;
32'b000000000000000000000000000001xx:y=5'b00010;
32'b00000000000000000000000000001xxx:y=5'b00011;
32'b0000000000000000000000000001xxxx:y=5'b00100;
32'b000000000000000000000000001xxxxx:y=5'b00101;
32'b00000000000000000000000001xxxxxx:y=5'b00110;
32'b0000000000000000000000001xxxxxxx:y=5'b00111;
32'b000000000000000000000001xxxxxxxx:y=5'b01000;
32'b00000000000000000000001xxxxxxxxx:y=5'b01001;
32'b0000000000000000000001xxxxxxxxxx:y=5'b01010;
32'b000000000000000000001xxxxxxxxxxx:y=5'b01011;
32'b00000000000000000001xxxxxxxxxxxx:y=5'b01100;
32'b0000000000000000001xxxxxxxxxxxxx:y=5'b01101;
32'b000000000000000001xxxxxxxxxxxxxx:y=5'b01110;
32'b00000000000000001xxxxxxxxxxxxxxx:y=5'b01111;
32'b0000000000000001xxxxxxxxxxxxxxxx:y=5'b10000;
32'b000000000000001xxxxxxxxxxxxxxxxx:y=5'b10001;
32'b00000000000001xxxxxxxxxxxxxxxxxx:y=5'b10010;
32'b0000000000001xxxxxxxxxxxxxxxxxxx:y=5'b10011;
32'b000000000001xxxxxxxxxxxxxxxxxxxx:y=5'b10100;
32'b00000000001xxxxxxxxxxxxxxxxxxxxx:y=5'b10101;
32'b0000000001xxxxxxxxxxxxxxxxxxxxxx:y=5'b10110;
32'b000000001xxxxxxxxxxxxxxxxxxxxxxx:y=5'b10111;
32'b00000001xxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11000;
32'b0000001xxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11001;
32'b000001xxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11010;
32'b00001xxxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11011;
32'b0001xxxxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11100;
32'b001xxxxxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11101;
32'b01xxxxxxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11110;
32'b1xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx:y=5'b11111;
default:y=5'bzzzzz;
endcase
end
endmodule
