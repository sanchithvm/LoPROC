`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer: Sanchith V M
//
// Create Date:    17:48:59 07/02/2022
// Design Name:
// Module Name:    loproc_defines
// Project Name: 	LoPROC v1.1
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`define DATA_WIDTH            32
`define INSTRUCTION_WIDTH     32
`define REG_BANK_DEPTH        32
`define REG_BANK_ADDR_WIDTH   5
`define DATA_LOG2             5
`define POWER_MODES           4
`define POWER_MODES_LOG2      2  
